entity main is
port(
end entity;
