LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_ARITH.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;

LIBRARY altera_mf;
USE altera_mf.all;

entity text_setter is
    PORT
    (
        character_address     :    OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
        pixel_row, pixel_col    :    IN STD_LOGIC_VECTOR (9 DOWNTO 4);
        clock                               :     IN STD_LOGIC ;
        rom_mux_output        :    OUT STD_LOGIC
    );
end text_setter;

architecture behave of text_setter is
begin

    process (pixel_col) 
    begin
        if(pixel_row= "00010") then
            if (pixel_col ="00010") then
                character_address <= "000110"; --F
            elsif (pixel_col ="00011") then
                character_address <= "001100"; --L
            elsif (pixel_col ="00100") then
                character_address <= "000001"; --A
            elsif (pixel_col ="00101") then
                character_address <= "010000"; --P
            elsif (pixel_col ="00111") then
                character_address <= "010000"; --P
            elsif (pixel_col ="01000") then
                character_address <= "000001"; --Y
            else
                character_address <= "100000";
            end if;
        else 
            character_address <= "100000";
        end if;
    end process;

end architecture;
